module controlUnit (
    
);
mainDeco mainDeco_1 (

);
aluDeco aluDeco_1(

);
endmodule